library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

entity INSTRUCTION_EXECUTE is
  Port ( 
        PC1: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ALUSRC: IN STD_LOGIC;
        RD1, RD2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        EXT_IMM: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        SA: IN STD_LOGIC;
        FUNCT: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        ALUOP:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        BRANCH_ADDRESS: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        ZERO: OUT STD_LOGIC;
        ALURES: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) 
  );
end INSTRUCTION_EXECUTE;

architecture Behavioral of INSTRUCTION_EXECUTE is
COMPONENT ALU IS
    Port (
        OP1, OP2:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        SA: IN STD_LOGIC;
        CONTROL: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
        ZERO:OUT STD_LOGIC;
        RES: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) 
    );
END COMPONENT;
SIGNAL SRC: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL CONTROL: STD_LOGIC_VECTOR(5 DOWNTO 0);
begin

CONTROL<=ALUOP & FUNCT;
SRC<=RD2 WHEN ALUSRC='0' ELSE EXT_IMM;

ALU1:ALU PORT MAP(
 OP1=>RD1,
 OP2=>SRC, 
 SA=>SA,
 CONTROL => CONTROL, ZERO=>ZERO, RES=>ALURES);
BRANCH_ADDRESS<=PC1+EXT_IMM;


end Behavioral;
