library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity MEMORY_UNIT is
    Port ( 
            CLK, EN: IN STD_LOGIC;
            MEMWRITE: IN STD_LOGIC;
            RD2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            ALURES_IN:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            ALURES_OUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            MEMDATA: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
end MEMORY_UNIT;

architecture Behavioral of MEMORY_UNIT is

TYPE MEMORY IS ARRAY(0 TO 255) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL MEM: MEMORY := (OTHERS=>X"0000");
begin

PROCESS(CLK, MEMWRITE, ALURES_IN) IS
BEGIN

IF RISING_EDGE(CLK) THEN
    IF MEMWRITE='1' AND EN='1' THEN 
    MEM(CONV_INTEGER(ALURES_IN))<=RD2;
    END IF;
END IF;


END PROCESS;
MEMDATA<=MEM(TO_INTEGER(UNSIGNED(ALURES_IN)));
ALURES_OUT<=ALURES_IN;


end Behavioral;
