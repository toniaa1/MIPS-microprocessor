library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
entity INSTRUCTION_FETCH is
 Port (
    CLK: IN STD_LOGIC;
--    RST: IN STD_LOGIC
    EN: IN STD_LOGIC;
    JUMP, PC_SRC:IN STD_LOGIC;
    JUMP_ADDR:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    BRANCH_ADDR: IN STD_LOGIC_VECTOR(15 downto 0);
    INSTR_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    INSTR1: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    PC1: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
    
end INSTRUCTION_FETCH;

architecture Behavioral of INSTRUCTION_FETCH is
TYPE INSTR_MEM IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL INSTRUCTION_MEMORY: INSTR_MEM:=(
X"208A",
X"2205",
X"2183",

X"0D40",
X"0E47",
X"10D1",

X"0E64",
X"0B65",
X"0F76",

X"36FF",
X"16D6",
X"9404",
X"012A",
X"01B3",
X"1130",
X"7000",
X"5C00",
X"BC02",
X"2481",
X"D412",
X"E000",
OTHERS=>X"0000");
SIGNAL PC:STD_LOGIC_VECTOR(15 DOWNTO 0):=(OTHERS=>'0');
SIGNAL PC_AUX, NEXT_ADDR, AUXSGN:STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ADDRESS:STD_LOGIC_VECTOR(15 DOWNTO 0);
begin

PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
--    IF RST='1' THEN
--        pc<=x"0000";
        IF EN='1' THEN
            PC<=NEXT_ADDR;
        END IF;
--    END IF;
END IF;
END PROCESS;

ADDRESS<=PC;

INSTR_OUT<=INSTRUCTION_MEMORY(to_integer(unsigned(ADDRESS)));
INSTR1<=INSTRUCTION_MEMORY(to_integer(unsigned(ADDRESS+1)));

PC_AUX<=PC+1;
PC1<=PC_AUX;

AUXSGN<=BRANCH_ADDR WHEN PC_SRC='1' ELSE PC_AUX;
NEXT_ADDR<=JUMP_ADDR WHEN JUMP='1' ELSE AUXSGN;


end Behavioral;
