library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


entity MIPS is
 port (
 clk : in std_logic;
 btn : in std_logic_vector(4 downto 0);
 sw : in std_logic_vector(15 downto 0);
 led : out std_logic_vector(15 downto 0);
 an : out std_logic_vector(3 downto 0);
 cat : out std_logic_vector(6 downto 0)
 );
end MIPS;

architecture Behavioral of MIPS is

COMPONENT INSTRUCTION_EXECUTE is
  Port ( 
        PC1: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ALUSRC: IN STD_LOGIC;
        RD1, RD2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        EXT_IMM: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        SA: IN STD_LOGIC;
        FUNCT: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        ALUOP:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        BRANCH_ADDRESS: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        ZERO: OUT STD_LOGIC;
        ALURES: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) 
  );
end COMPONENT;

COMPONENT INSTRUCTION_DECODE is
  Port ( CLK: IN STD_LOGIC;
         EN: IN STD_LOGIC;
         REG_WRITE: IN STD_LOGIC;
         REGDst:IN STD_LOGIC;
         EXTop:IN STD_LOGIC;
         INSTR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
         WD:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
         RD1: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
         RD2: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
         FUNC: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
         SA:OUT STD_LOGIC;      
         EXT_IMM:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
         
end COMPONENT;

COMPONENT INSTRUCTION_FETCH is
 Port (
    CLK: IN STD_LOGIC;
--    RST: IN STD_LOGIC,
    EN: IN STD_LOGIC;
    JUMP, PC_SRC:IN STD_LOGIC;
    JUMP_ADDR:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    BRANCH_ADDR: IN STD_LOGIC_VECTOR(15 downto 0);
    INSTR_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    INSTR1: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    PC1: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
    
end COMPONENT;

COMPONENT MAIN_CONTROL is
Port ( 
        INSTR: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        ALUOP: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        REGDST, EXTOP, ALUSRC, BRANCH, JUMP, MEMWRITE, MEMTOREG, REGWRITE: OUT STD_LOGIC
);
end COMPONENT;

COMPONENT MEMORY_UNIT is
    Port ( 
            CLK, EN: IN STD_LOGIC;
            MEMWRITE: IN STD_LOGIC;
            RD2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            ALURES_IN:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            ALURES_OUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            MEMDATA: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
end COMPONENT;

COMPONENT SSD_DRIVER is
  Port (
    CLK: IN STD_LOGIC;
    NUM1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    NUM2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    NUM3: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    NUM4: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    an : out std_logic_vector(3 downto 0);
    cat : out std_logic_vector(6 downto 0));
END COMPONENT;

COMPONENT MPG is
  Port (BTN: IN STD_LOGIC;
         CLK:IN STD_LOGIC;
         BTNO:OUT STD_LOGIC);
END COMPONENT;

SIGNAL INSTR, INSTR1:STD_LOGIC_VECTOR(15 DOWNTO 0); 
SIGNAL REGDST, EXTOP, ALUSRC, BRANCH, JUMP, MEMWRITE, MEMTOREG, REGWRITE: STD_LOGIC; 
SIGNAL ZERO,PCSRC, BTNO: STD_LOGIC;
SIGNAL ALUOP: STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL JUMP_ADDR, BRANCH_ADDRESS, PC2, ALURES, ALURES1: STD_LOGIC_VECTOR(15 DOWNTO 0);
signal PC1,WD:STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RD1,RD2:STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FUNC: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL SA:STD_LOGIC;
SIGNAL EXT_IMM, MEMDATA:STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL NUM1, NUM2, NUM3, NUM4: STD_LOGIC_VECTOR(3 DOWNTO 0);

begin

IFETCH: INSTRUCTION_FETCH 
 Port MAP(
    CLK=>CLK,
--    RST=>SW(0),
    EN=>BTNO,
    JUMP=>JUMP, 
    PC_SRC=>PCSRC,
    JUMP_ADDR=>JUMP_ADDR,
    BRANCH_ADDR=>BRANCH_ADDRESS,
    INSTR_OUT=>INSTR,
    INSTR1=>INSTR1,
    PC1=>PC1);

ID:INSTRUCTION_DECODE 
  Port MAP ( CLK=>CLK,
            EN=>'1',
         REG_WRITE=>REGWRITE,
         REGDst=>REGDST,
         EXTop=>EXTOP,
         INSTR=>INSTR,
         WD=>WD,
         RD1=>RD1,
         RD2=>RD2,
         FUNC=>FUNC,
         SA=>SA,      
         EXT_IMM=>EXT_IMM);

MC:MAIN_CONTROL 
Port MAP( 
        INSTR=>INSTR(15 DOWNTO 13),
        ALUOP=>ALUOP,
        REGDST=>REGDST, 
        EXTOP=>EXTOP, 
        ALUSRC=>ALUSRC, 
        BRANCH=>BRANCH,
        JUMP=>JUMP, 
        MEMWRITE=>MEMWRITE, 
        MEMTOREG=>MEMTOREG, 
        REGWRITE=>REGWRITE);

IE: INSTRUCTION_EXECUTE PORT MAP ( 
        PC1=>PC1,
        ALUSRC=>ALUSRC,
        RD1=>RD1,
        RD2=>RD2,
        EXT_IMM=>EXT_IMM,
        SA=>SA,
        FUNCT=>FUNC,
        ALUOP=>ALUOP,
        BRANCH_ADDRESS=>BRANCH_ADDRESS,
        ZERO=>ZERO,
        ALURES=>ALURES);

MU:MEMORY_UNIT Port MAP( 
            CLK=>CLK, 
            EN=>BTNO,
            MEMWRITE=>MEMWRITE,
            RD2=>RD2,
            ALURES_IN=>ALURES,
            ALURES_OUT=>ALURES1,
            MEMDATA=>MEMDATA);

MPG1: MPG PORT MAP(BTN=>BTN(0), CLK=>CLK, BTNO=>BTNO);
SSD: SSD_DRIVER PORT MAP(CLK=>CLK, 
                         NUM1=>NUM1, 
                         NUM2=>NUM2, 
                         NUM3=>NUM3, 
                         NUM4=>NUM4, 
                         AN=>AN, 
                         CAT=>CAT);




WD <= MemData when MemtoReg = '1' else ALURes1;
PCSRC<=ZERO AND BRANCH;
JUMP_ADDR<=PC1(15 DOWNTO 13) & INSTR(12 DOWNTO 0);

PROCESS(SW, INSTR, INSTR1, RD1, RD2, EXT_IMM, ALURES, MEMDATA, WD) IS 
BEGIN

CASE(SW (7 DOWNTO 5)) IS
WHEN "000"=>
    NUM1<=INSTR(15 DOWNTO 12);
    NUM2<=INSTR(11 DOWNTO 8);
    NUM3<=INSTR(7 DOWNTO 4);
    NUM4<=INSTR(3 DOWNTO 0);
WHEN "001"=>
    NUM1<=INSTR1(15 DOWNTO 12);
    NUM2<=INSTR1(11 DOWNTO 8);
    NUM3<=INSTR1(7 DOWNTO 4);
    NUM4<=INSTR1(3 DOWNTO 0);
WHEN "010"=>
    NUM1<=RD1(15 DOWNTO 12);
    NUM2<=RD1(11 DOWNTO 8);
    NUM3<=RD1(7 DOWNTO 4);
    NUM4<=RD1(3 DOWNTO 0);
WHEN "011"=>
    NUM1<=RD2(15 DOWNTO 12);
    NUM2<=RD2(11 DOWNTO 8);
    NUM3<=RD2(7 DOWNTO 4);
    NUM4<=RD2(3 DOWNTO 0);
WHEN "100"=>
    NUM1<=EXT_IMM(15 DOWNTO 12);
    NUM2<=EXT_IMM(11 DOWNTO 8);
    NUM3<=EXT_IMM(7 DOWNTO 4);
    NUM4<=EXT_IMM(3 DOWNTO 0);
WHEN "101"=>
    NUM1<=ALURES(15 DOWNTO 12);
    NUM2<=ALURES(11 DOWNTO 8);
    NUM3<=ALURES(7 DOWNTO 4);
    NUM4<=ALURES(3 DOWNTO 0);
WHEN "110"=>
    NUM1<=MEMDATA(15 DOWNTO 12);
    NUM2<=MEMDATA(11 DOWNTO 8);
    NUM3<=MEMDATA(7 DOWNTO 4);
    NUM4<=MEMDATA(3 DOWNTO 0);
WHEN "111"=>
    NUM1<=WD(15 DOWNTO 12);
    NUM2<=WD(11 DOWNTO 8);
    NUM3<=WD(7 DOWNTO 4);
    NUM4<=WD(3 DOWNTO 0);
END CASE;

    LED(0)<=ALUSRC;
    LED(1)<=MEMWRITE;
    LED(2)<=MEMTOREG;
    LED(3)<=REGWRITE;
    LED(4)<=JUMP;
    LED(5)<=BRANCH;
    LED(6)<=EXTOP;
    LED(7)<=REGDST;
    
    led(8)<=btno;
    
    LED(10)<=ALUOP(0);
    LED(11)<=ALUOP(1);
    LED(12)<=ALUOP(2);
    LED(15)<=ZERO;
end process;

end Behavioral;
