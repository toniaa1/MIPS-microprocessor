library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

entity MPG is
  Port (BTN: IN STD_LOGIC;
         CLK:IN STD_LOGIC;
         BTNO:OUT STD_LOGIC);
end MPG;

architecture Behavioral of MPG is

SIGNAL D1, D2, D3: STD_LOGIC;
SIGNAL COUNT:STD_LOGIC_VECTOR (15 DOWNTO 0);
begin

PROCESS(CLK) IS
BEGIN
IF RISING_EDGE(CLK) THEN
    COUNT<=COUNT+1;
END IF;
END PROCESS;



PROCESS(COUNT, CLK) IS
BEGIN

IF RISING_EDGE(CLK) THEN
IF COUNT =X"FFFF" THEN
    D1<=BTN;
END IF;
END IF;   
END PROCESS;

PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
    D2<=D1;
    D3<=D2;
END IF;
END PROCESS;


BTNO<=NOT D3 AND D2;


end Behavioral;
